module main

fn main() {
	println('Hello World!')
	nums := []int{len: 10, init: it}
	println(nums)
	dbls := nums.map(it * 2)
	println(dbls)
	sqrs := nums.map(it * it)
	println(sqrs)
}
